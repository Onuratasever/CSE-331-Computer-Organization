module my_or_32bit( 
							output [31:0]out,
							input [31:0]a,
							input [31:0]b

						); 


or or1(out[0],a[0],b[0]);
or or2(out[1],a[1],b[1]);
or or3(out[2],a[2],b[2]);
or or4(out[3],a[3],b[3]);
or or5(out[4],a[4],b[4]);
or or6(out[5],a[5],b[5]);
or or7(out[6],a[6],b[6]);
or or8(out[7],a[7],b[7]);
or or9(out[8],a[8],b[8]);
or or10(out[9],a[9],b[9]);
or or11(out[10],a[10],b[10]);
or or12(out[11],a[11],b[11]);
or or13(out[12],a[12],b[12]);
or or14(out[13],a[13],b[13]);
or or15(out[14],a[14],b[14]);
or or16(out[15],a[15],b[15]);
or or17(out[16],a[16],b[16]);
or or18(out[17],a[17],b[17]);
or or19(out[18],a[18],b[18]);
or or20(out[19],a[19],b[19]);
or or21(out[20],a[20],b[20]);
or or22(out[21],a[21],b[21]);
or or23(out[22],a[22],b[22]);
or or24(out[23],a[23],b[23]);
or or25(out[24],a[24],b[24]);
or or26(out[25],a[25],b[25]);
or or27(out[26],a[26],b[26]);
or or28(out[27],a[27],b[27]);
or or29(out[28],a[28],b[28]);
or or30(out[29],a[29],b[29]);
or or31(out[30],a[30],b[30]);
or or32(out[31],a[31],b[31]);

endmodule
