module extend_32bit( //
	output [31:1] out,
	input a,
	input b
); 


or or2(out[1],a,b);
or or3(out[2],a,b);
or or4(out[3],a,b);
or or5(out[4],a,b);
or or6(out[5],a,b);
or or7(out[6],a,b);
or or8(out[7],a,b);
or or9(out[8],a,b);
or or10(out[9],a,b);
or or11(out[10],a,b);
or or12(out[11],a,b);
or or13(out[12],a,b);
or or14(out[13],a,b);
or or15(out[14],a,b);
or or16(out[15],a,b);
or or17(out[16],a,b);
or or18(out[17],a,b);
or or19(out[18],a,b);
or or20(out[19],a,b);
or or21(out[20],a,b);
or or22(out[21],a,b);
or or23(out[22],a,b);
or or24(out[23],a,b);
or or25(out[24],a,b);
or or26(out[25],a,b);
or or27(out[26],a,b);
or or28(out[27],a,b);
or or29(out[28],a,b);
or or30(out[29],a,b);
or or31(out[30],a,b);
or or32(out[31],a,b);

endmodule
